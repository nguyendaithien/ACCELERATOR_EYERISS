module PE #(parameter DATA_IN_WIDTH = 8, DATA_OUT_WIDTH = 16)(
		clk,
		rst_n,
		ifm,
		wgt,
		psum_in,
    psum_out,
		set_wgt,
		
